//`define RISKV_DEBUG 0
